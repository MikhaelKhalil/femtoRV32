`timescale 1ns / 1ps

module InstMem(
	input [7:0] addr,
	output [31:0] data_out
    );

    // reg [31:0] mem [0:255];  // change into 8 bits when using at byte-addressable
	reg [31:0] mem [0:255];
	assign data_out = mem[addr];

	initial begin
        /* COMPREHENSIVE TEST PROGRAM */
        mem[0] = 32'b00010010001101000101000010110111;      // LUI   x1, 0x12345    # 0x12345000
        mem[4] = 32'b00000000000000010000000100010111;      // AUIPC x2, 0x10       # 0x10000
        mem[8] = 32'b00000000010100001000000110010011;      // ADDI  x3, x1, 5      # 305418245
        mem[12] = 32'b00000000101000011010001000010011;      // SLTI  x4, x3, 10    # 0
        mem[16] = 32'b00000000100100011011001010010011;      // SLTIU x5, x3, 9     # 0
        mem[20] = 32'b00000000100000011100001100010011;      // XORI  x6, x3, 8     # 305418253
        mem[24] = 32'b00000000011100011110001110010011;      // ORI   x7, x3, 7     # 305418247
        mem[28] = 32'b00000000001100011111010000010011;      // ANDI  x8, x3, 3     # 1
        mem[32] = 32'b00000000001000011001010010010011;      // SLLI  x9, x3, 2     # 1221672980
        mem[36] = 32'b00000000000100011101010100010011;      // SRLI  x10, x3, 1    # 152709122
        mem[40] = 32'b01000000000100011101010110010011;     // SRAI  x11, x3, 1     # 152709122
        mem[44] = 32'b00000000000100011000011000110011;     // ADD   x12, x3, x1    # 610836485
        mem[48] = 32'b01000000000100011000011010110011;     // SUB   x13, x3, x1    # 5
        mem[52] = 32'b00000000110100011001011100110011;     // SLL   x14, x3, x13   # 9773383840 => clipped into => 1183449248
        mem[56] = 32'b00000000001100001010011110110011;     // SLT   x15, x1, x3    # 1
        mem[60] = 32'b00000000000100011011100000110011;     // SLTU  x16, x3, x1    # 0
        mem[64] = 32'b00000000000100011100100010110011;     // XOR   x17, x3, x1    # 5
        mem[68] = 32'b00000000110100011101100100110011;     // SRL   x18, x3, x13   # 9544320
        mem[72] = 32'b01000000110100011101100110110011;     // SRA   x19, x3, x13   # 9544320
        mem[76] = 32'b00000000000100011110101000110011;     // OR    x20, x3, x1    # 305418245
        mem[80] = 32'b00000000000100011111101010110011;     // AND   x21, x3, x1    # 305418240
        mem[84] = 32'b00000000001100000010000000100011;     // SW    x3, 0(x0)      # mem[3:0] changed
        mem[88] = 32'b00000000001100000001001000100011;     // SH    x3, 4(x0)      # mem[5:4] changed 
        mem[92] = 32'b00000000001100000000001100100011;     // SB    x3, 6(x0)      # mem[6] changed
        mem[96] = 32'b00000000000000000010101100000011;     // LW    x22, 0(x0)     # 305418245
        mem[100] = 32'b00000000010000000001101110000011;     // LH    x23, 4(x0)    # 
        mem[104] = 32'b00000000011000000000110000000011;     // LB    x24, 6(x0)    # 5
        mem[108] = 32'b00000000010000000101110010000011;     // LHU   x25, 4(x0)    # 
        mem[112] = 32'b00000000011000000100110100000011;     // LBU   x26, 6(x0)    # 5
        mem[116] = 32'b00000000010100000000110110010011;     // ADDI  x27, x0, 5    # 5
        mem[120] = 32'b00000000101000000000111000010011;     // ADDI  x28, x0, 10   # 10
        mem[124] = 32'b00000001110011011000010001100011;     // BEQ   x27, x28, skip_beq                # not taken
        mem[128] = 32'b00000000000100000000111010010011;     // ADDI  x29, x0, 1                        # 1
        mem[132] = 32'b00000001110011011001010001100011;     // skip_beq: BNE   x27, x28, after_bne     # taken => 140
        mem[136] = 32'b00000000001000000000111010010011;     // ADDI  x29, x0, 2
        mem[140] = 32'b00000001110011011100010001100011;     // after_bne: BLT   x27, x28, after_blt    # 5 < 10 => taken => 148
        mem[144] = 32'b00000000001100000000111100010011;     // ADDI  x30, x0, 3
        mem[148] = 32'b00000001101111100101010001100011;     // after_blt: BGE   x28, x27, after_bge    # 10 > 5 => taken => 156
        mem[152] = 32'b00000000010000000000111100010011;     // ADDI  x30, x0, 4
        mem[156] = 32'b00000001101111100110010001100011;     // after_bge: BLTU  x28, x27, after_bltu   # 10 !< 5 => not taken
        mem[160] = 32'b00000000010100000000111100010011;     // ADDI  x30, x0, 5                        # 5
        mem[164] = 32'b00000001110011011111010001100011;     // after_bltu: BGEU  x27, x28, after_bgeu  # 5 !> 10 => not taken
        mem[168] = 32'b00000000011000000000111100010011;     // ADDI  x30, x0, 6                        # 6
        mem[172] = 32'b00000000100000000000111111101111;     // after_bgeu: JAL   x31, jal_target       # PC => 180, x31 => 176
        mem[176] = 32'b00000110001100000000001010010011;     // ADDI  x5, x0, 99
        mem[180] = 32'b00000010101000000000001100010011;     // jal_target: ADDI  x6, x0, 42            # 42
        // mem[184] = 32'b00000000000011111000010101100111;     // JALR  x10, x31, 0                       # PC => 176, x10 => 188
        // mem[184] = 32'b00000000000000000001000000001111;     // FENCE.I
        mem[184] = 32'b00000000000000000000000001110011;     // ECALL
        // mem[184] = 32'b00000000000100000000000001110011;     // EBREAK
        mem[188] = 32'b00000000000011111000010101100111;        // JALR  x10, x31, 0                       # PC => 176, x10 => 188
	end

endmodule
